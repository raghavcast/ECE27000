(* blackbox *)
module hangman (
  input logic hz100, reset, flash,
  input logic [5:0] hex,
  output logic [6:0] ctrdisp,
  output logic [27:0] letterdisp,
  output logic win, lose
);

// This file is INTENTIONALLY empty!
// Do not enter any code here! - NM

endmodule